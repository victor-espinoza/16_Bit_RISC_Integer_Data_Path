`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
// Author:         Victor Espinoza
// Partner:        Edward Mares
// Email:          victor.alfonso94@gmail.com
// 
// Create Date:    19:42:15 10/12/2013 
// Module Name:    ad_mux 
// File Name:      ad_mux.v
// 
// Description:    This multiplexer mudule is used to select what data input are to 
//                 be assigned to the ad_out output and driven to the seven segment
//                 display. The value of the ad_out is chosen based on the seg_sel
//                 input that was generated by our led_controller module.
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ad_mux(seg_sel, ad_high, ad_low, d_high, d_low, ad_out);

   //Inputs
   input          [1:0] seg_sel;
   input          [3:0] ad_high, ad_low, d_high, d_low;
   
   //Ouput
   output         [3:0] ad_out;
   reg            [3:0] ad_out;
   
   always @(seg_sel or ad_high or ad_low or d_high or d_low)   
      case (seg_sel)      
         2'b00  :      ad_out =  d_low;    //annode 0
         2'b01  :      ad_out =  d_high;   //annode 1
         2'b10  :      ad_out =  ad_low;   //annode 2
         2'b11  :      ad_out =  ad_high;  //annode 3
         default:    ad_out =  1'bx;  //default output   
      endcase      
endmodule
